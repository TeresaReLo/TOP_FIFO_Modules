module fv_top_module#(

);



/////// Assumptionss//////////////////////
  

/////// Assertions //////////////////////
   
   
/////// Cover properties/////////////////
        


endmodule


bind top_module fv_top_module fv_top_module_inst(.*);
