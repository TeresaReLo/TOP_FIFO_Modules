/* 
	=========================================================================================
	Module name	: funct_generator LUT
	Author		: Ana Godoy
	Email		: ana.gm@circuify.com
	Filename	: funct_generator_lut.sv
	Type		: SystemVerilog Module
	
	Description	:LUT
	-----------------------------------------------------------------------------------------
		clocks	: clk

	-----------------------------------------------------------------------------------------
	Version		: 1.0
	Date		: Jun 2024
	-----------------------------------------------------------------------------------------
*/

module funct_generator_lut #(
		parameter DATA_WIDTH= 32,
		parameter ADDR_WIDTH= 8,
		parameter TXT_FILE= "sin.txt"
)(
		//Inputs
		input  logic                  clk,		
		input  logic [ADDR_WIDTH-1:0] read_addr_i,
		//Outputs
		output logic signed [DATA_WIDTH-1 : 0] read_data_o
);

// signal declaration
	reg [DATA_WIDTH-1:0] lut_structure [2**ADDR_WIDTH-1:0]; 
/*
initial begin  //load hexadecimal data in txt
		//$readmemh(TXT_FILE, lut_structure);

                //sine
                if(TXT_FILE == 1) begin
                    lut_structure[0]   = 32'h00000000;
                    lut_structure[1]   = 32'h00645A1C;
                    lut_structure[2]   = 32'h00C91D14;
                    lut_structure[3]   = 32'h012D7731;
                    lut_structure[4]   = 32'h01916872;
                    lut_structure[5]   = 32'h01F559B3;
                    lut_structure[6]   = 32'h0258E219;
                    lut_structure[7]   = 32'h02BC6A7E;
                    lut_structure[8]   = 32'h031F212D;
                    lut_structure[9]   = 32'h03816F00;
                    lut_structure[10]  = 32'h03E353F7;
                    lut_structure[11]  = 32'h04446738;
                    lut_structure[12]  = 32'h04A5119C;
                    lut_structure[13]  = 32'h0504EA4A;
                    lut_structure[14]  = 32'h0563F141;
                    lut_structure[15]  = 32'h05C22680;
                    lut_structure[16]  = 32'h061F8A09;
                    lut_structure[17]  = 32'h067BB2FE;
                    lut_structure[18]  = 32'h06D77318;
                    lut_structure[19]  = 32'h07318FC5;
                    lut_structure[20]  = 32'h078ADAB9;
                    lut_structure[21]  = 32'h07E2EB1C;
                    lut_structure[22]  = 32'h0839C0EB;
                    lut_structure[23]  = 32'h088F5C28;
                    lut_structure[24]  = 32'h08E3BCD3;
                    lut_structure[25]  = 32'h09367A0F;
                    lut_structure[26]  = 32'h0987FCB9;
                    lut_structure[27]  = 32'h09D7DBF4;
                    lut_structure[28]  = 32'h0A26809D;
                    lut_structure[29]  = 32'h0A7381D7;
                    lut_structure[30]  = 32'h0ABEDFA4;
                    lut_structure[31]  = 32'h0B083126;
                    lut_structure[32]  = 32'h0B504816;
                    lut_structure[33]  = 32'h0B9652BD;
                    lut_structure[34]  = 32'h0BDB22D0;
                    lut_structure[35]  = 32'h0C1D7DBF;
                    lut_structure[36]  = 32'h0C5E353F;
                    lut_structure[37]  = 32'h0C9CE075;
                    lut_structure[38]  = 32'h0CD9E83E;
                    lut_structure[39]  = 32'h0D14E3BC;
                    lut_structure[40]  = 32'h0D4DD2F1;
                    lut_structure[41]  = 32'h0D84B5DC;
                    lut_structure[42]  = 32'h0DB923A2;
                    lut_structure[43]  = 32'h0DEBEDFA;
                    lut_structure[44]  = 32'h0E1C432C;
                    lut_structure[45]  = 32'h0E4A8C15;
                    lut_structure[46]  = 32'h0E76C8B4;
                    lut_structure[47]  = 32'h0EA0902D;
                    lut_structure[48]  = 32'h0EC84B5D;
                    lut_structure[49]  = 32'h0EED9168;
                    lut_structure[50]  = 32'h0F10624D;
                    lut_structure[51]  = 32'h0F3126E9;
                    lut_structure[52]  = 32'h0F4F765F;
                    lut_structure[53]  = 32'h0F6BB98C;
                    lut_structure[54]  = 32'h0F851EB8;
                    lut_structure[55]  = 32'h0F9C779A;
                    lut_structure[56]  = 32'h0FB15B57;
                    lut_structure[57]  = 32'h0FC3C9EE;
                    lut_structure[58]  = 32'h0FD3C361;
                    lut_structure[59]  = 32'h0FE147AE;
                    lut_structure[60]  = 32'h0FEC56D5;
                    lut_structure[61]  = 32'h0FF4F0D8;
                    lut_structure[62]  = 32'h0FFB15B5;
                    lut_structure[63]  = 32'h0FFEC56D;
                    lut_structure[64]  = 32'h10000000;
                    lut_structure[65]  = 32'h0FFEC56D;
                    lut_structure[66]  = 32'h0FFB15B5;
                    lut_structure[67]  = 32'h0FF4F0D8;
                    lut_structure[68]  = 32'h0FEC56D5;
                    lut_structure[69]  = 32'h0FE147AE;
                    lut_structure[70]  = 32'h0FD3C361;
                    lut_structure[71]  = 32'h0FC3C9EE;
                    lut_structure[72]  = 32'h0FB15B57;
                    lut_structure[73]  = 32'h0F9C779A;
                    lut_structure[74]  = 32'h0F851EB8;
                    lut_structure[75]  = 32'h0F6BB98C;
                    lut_structure[76]  = 32'h0F4F765F;
                    lut_structure[77]  = 32'h0F3126E9;
                    lut_structure[78]  = 32'h0F10624D;
                    lut_structure[79]  = 32'h0EED9168;
                    lut_structure[80]  = 32'h0EC84B5D;
                    lut_structure[81]  = 32'h0EA0902D;
                    lut_structure[82]  = 32'h0E76C8B4;
                    lut_structure[83]  = 32'h0E4A8C15;
                    lut_structure[84]  = 32'h0E1C432C;
                    lut_structure[85]  = 32'h0DEBEDFA;
                    lut_structure[86]  = 32'h0DB923A2;
                    lut_structure[87]  = 32'h0D84B5DC;
                    lut_structure[88]  = 32'h0D4DD2F1;
                    lut_structure[89]  = 32'h0D14E3BC;
                    lut_structure[90]  = 32'h0CD9E83E;
                    lut_structure[91]  = 32'h0C9CE075;
                    lut_structure[92]  = 32'h0C5E353F;
                    lut_structure[93]  = 32'h0C1D7DBF;
                    lut_structure[94]  = 32'h0BDB22D0;
                    lut_structure[95]  = 32'h0B9652BD;
                    lut_structure[96]  = 32'h0B504816;
                    lut_structure[97]  = 32'h0B083126;
                    lut_structure[98]  = 32'h0ABEDFA4;
                    lut_structure[99]  = 32'h0A7381D7;
                    lut_structure[100] = 32'h0A26809D;
                    lut_structure[101] = 32'h09D7DBF4;
                    lut_structure[102] = 32'h0987FCB9;
                    lut_structure[103] = 32'h09367A0F;
                    lut_structure[104] = 32'h08E3BCD3;
                    lut_structure[105] = 32'h088F5C28;
                    lut_structure[106] = 32'h0839C0EB;
                    lut_structure[107] = 32'h07E2EB1C;
                    lut_structure[108] = 32'h078ADAB9;
                    lut_structure[109] = 32'h07318FC5;
                    lut_structure[110] = 32'h06D77318;
                    lut_structure[111] = 32'h067BB2FE;
                    lut_structure[112] = 32'h061F8A09;
                    lut_structure[113] = 32'h05C22680;
                    lut_structure[114] = 32'h0563F141;
                    lut_structure[115] = 32'h0504EA4A;
                    lut_structure[116] = 32'h04A5119C;
                    lut_structure[117] = 32'h04446738;
                    lut_structure[118] = 32'h03E353F7;
                    lut_structure[119] = 32'h03816F00;
                    lut_structure[120] = 32'h031F212D;
                    lut_structure[121] = 32'h02BC6A7E;
                    lut_structure[122] = 32'h0258E219;
                    lut_structure[123] = 32'h01F559B3;
                    lut_structure[124] = 32'h01916872;
                    lut_structure[125] = 32'h012D7731;
                    lut_structure[126] = 32'h00C91D14;
                    lut_structure[127] = 32'h00645A1C;
                    lut_structure[128] = 32'h00000000;
                    lut_structure[129] = 32'hFF9BA5E4;
                    lut_structure[130] = 32'hFF36E2EC;
                    lut_structure[131] = 32'hFED288CF;
                    lut_structure[132] = 32'hFE6E978E;
                    lut_structure[133] = 32'hFE0AA64D;
                    lut_structure[134] = 32'hFDA71DE7;
                    lut_structure[135] = 32'hFD439582;
                    lut_structure[136] = 32'hFCE0DED3;
                    lut_structure[137] = 32'hFC7E91FF;
                    lut_structure[138] = 32'hFC1CAC09;
                    lut_structure[139] = 32'hFBBB98C8;
                    lut_structure[140] = 32'hFB5AEE64;
                    lut_structure[141] = 32'hFAFB15B6;
                    lut_structure[142] = 32'hFA9C0EBF;
                    lut_structure[143] = 32'hFA3DD980;
                    lut_structure[144] = 32'hF9E075F7;
                    lut_structure[145] = 32'hF9844D02;
                    lut_structure[146] = 32'hF9288CE8;
                    lut_structure[147] = 32'hF8CE703B;
                    lut_structure[148] = 32'hF8752547;
                    lut_structure[149] = 32'hF81D14E4;
                    lut_structure[150] = 32'hF7C63F15;
                    lut_structure[151] = 32'hF770A3D8;
                    lut_structure[152] = 32'hF71C432D;
                    lut_structure[153] = 32'hF6C985F1;
                    lut_structure[154] = 32'hF6780347;
                    lut_structure[155] = 32'hF628240C;
                    lut_structure[156] = 32'hF5D97F63;
                    lut_structure[157] = 32'hF58C7E29;
                    lut_structure[158] = 32'hF541205C;
                    lut_structure[159] = 32'hF4F7CEDA;
                    lut_structure[160] = 32'hF4AFB7EA;
                    lut_structure[161] = 32'hF469AD43;
                    lut_structure[162] = 32'hF424DD30;
                    lut_structure[163] = 32'hF3E28241;
                    lut_structure[164] = 32'hF3A1CAC1;
                    lut_structure[165] = 32'hF3631F8B;
                    lut_structure[166] = 32'hF32617C2;
                    lut_structure[167] = 32'hF2EB1C44;
                    lut_structure[168] = 32'hF2B22D0F;
                    lut_structure[169] = 32'hF27B4A24;
                    lut_structure[170] = 32'hF246DC5E;
                    lut_structure[171] = 32'hF2141206;
                    lut_structure[172] = 32'hF1E3BCD4;
                    lut_structure[173] = 32'hF1B573EB;
                    lut_structure[174] = 32'hF189374C;
                    lut_structure[175] = 32'hF15F6FD3;
                    lut_structure[176] = 32'hF137B4A3;
                    lut_structure[177] = 32'hF1126E98;
                    lut_structure[178] = 32'hF0EF9DB3;
                    lut_structure[179] = 32'hF0CED917;
                    lut_structure[180] = 32'hF0B089A1;
                    lut_structure[181] = 32'hF0944674;
                    lut_structure[182] = 32'hF07AE148;
                    lut_structure[183] = 32'hF0638866;
                    lut_structure[184] = 32'hF04EA4A9;
                    lut_structure[185] = 32'hF03C3612;
                    lut_structure[186] = 32'hF02C3C9F;
                    lut_structure[187] = 32'hF01EB852;
                    lut_structure[188] = 32'hF013A92B;
                    lut_structure[189] = 32'hF00B0F28;
                    lut_structure[190] = 32'hF004EA4B;
                    lut_structure[191] = 32'hF0013A93;
                    lut_structure[192] = 32'hF0000000;
                    lut_structure[193] = 32'hF0013A93;
                    lut_structure[194] = 32'hF004EA4B;
                    lut_structure[195] = 32'hF00B0F28;
                    lut_structure[196] = 32'hF013A92B;
                    lut_structure[197] = 32'hF01EB852;
                    lut_structure[198] = 32'hF02C3C9F;
                    lut_structure[199] = 32'hF03C3612;
                    lut_structure[200] = 32'hF04EA4A9;
                    lut_structure[201] = 32'hF0638866;
                    lut_structure[202] = 32'hF07AE148;
                    lut_structure[203] = 32'hF0944674;
                    lut_structure[204] = 32'hF0B089A1;
                    lut_structure[205] = 32'hF0CED917;
                    lut_structure[206] = 32'hF0EF9DB3;
                    lut_structure[207] = 32'hF1126E98;
                    lut_structure[208] = 32'hF137B4A3;
                    lut_structure[209] = 32'hF15F6FD3;
                    lut_structure[210] = 32'hF189374C;
                    lut_structure[211] = 32'hF1B573EB;
                    lut_structure[212] = 32'hF1E3BCD4;
                    lut_structure[213] = 32'hF2141206;
                    lut_structure[214] = 32'hF246DC5E;
                    lut_structure[215] = 32'hF27B4A24;
                    lut_structure[216] = 32'hF2B22D0F;
                    lut_structure[217] = 32'hF2EB1C44;
                    lut_structure[218] = 32'hF32617C2;
                    lut_structure[219] = 32'hF3631F8B;
                    lut_structure[220] = 32'hF3A1CAC1;
                    lut_structure[221] = 32'hF3E28241;
                    lut_structure[222] = 32'hF424DD30;
                    lut_structure[223] = 32'hF469AD43;
                    lut_structure[224] = 32'hF4AFB7EA;
                    lut_structure[225] = 32'hF4F7CEDA;
                    lut_structure[226] = 32'hF541205C;
                    lut_structure[227] = 32'hF58C7E29;
                    lut_structure[228] = 32'hF5D97F63;
                    lut_structure[229] = 32'hF628240C;
                    lut_structure[230] = 32'hF6780347;
                    lut_structure[231] = 32'hF6C985F1;
                    lut_structure[232] = 32'hF71C432D;
                    lut_structure[233] = 32'hF770A3D8;
                    lut_structure[234] = 32'hF7C63F15;
                    lut_structure[235] = 32'hF81D14E4;
                    lut_structure[236] = 32'hF8752547;
                    lut_structure[237] = 32'hF8CE703B;
                    lut_structure[238] = 32'hF9288CE8;
                    lut_structure[239] = 32'hF9844D02;
                    lut_structure[240] = 32'hF9E075F7;
                    lut_structure[241] = 32'hFA3DD980;
                    lut_structure[242] = 32'hFA9C0EBF;
                    lut_structure[243] = 32'hFAFB15B6;
                    lut_structure[244] = 32'hFB5AEE64;
                    lut_structure[245] = 32'hFBBB98C8;
                    lut_structure[246] = 32'hFC1CAC09;
                    lut_structure[247] = 32'hFC7E91FF;
                    lut_structure[248] = 32'hFCE0DED3;
                    lut_structure[249] = 32'hFD439582;
                    lut_structure[250] = 32'hFDA71DE7;
                    lut_structure[251] = 32'hFE0AA64D;
                    lut_structure[252] = 32'hFE6E978E;
                    lut_structure[253] = 32'hFED288CF;
                    lut_structure[254] = 32'hFF36E2EC;
                    lut_structure[255] = 32'hFF9BA5E4; 
                end
                //cosine
                else if(TXT_FILE == 2) begin
                    lut_structure[0]   = 32'h10000000;
                    lut_structure[1]   = 32'h0FFEC56D;
                    lut_structure[2]   = 32'h0FFB15B5;
                    lut_structure[3]   = 32'h0FF4F0D8;
                    lut_structure[4]   = 32'h0FEC56D5;
                    lut_structure[5]   = 32'h0FE147AE;
                    lut_structure[6]   = 32'h0FD3C361;
                    lut_structure[7]   = 32'h0FC3C9EE;
                    lut_structure[8]   = 32'h0FB15B57;
                    lut_structure[9]   = 32'h0F9C779A;
                    lut_structure[10]  = 32'h0F851EB8;
                    lut_structure[11]  = 32'h0F6BB98C;
                    lut_structure[12]  = 32'h0F4F765F;
                    lut_structure[13]  = 32'h0F3126E9;
                    lut_structure[14]  = 32'h0F10624D;
                    lut_structure[15]  = 32'h0EED9168;
                    lut_structure[16]  = 32'h0EC84B5D;
                    lut_structure[17]  = 32'h0EA0902D;
                    lut_structure[18]  = 32'h0E76C8B4;
                    lut_structure[19]  = 32'h0E4A8C15;
                    lut_structure[20]  = 32'h0E1C432C;
                    lut_structure[21]  = 32'h0DEBEDFA;
                    lut_structure[22]  = 32'h0DB923A2;
                    lut_structure[23]  = 32'h0D84B5DC;
                    lut_structure[24]  = 32'h0D4DD2F1;
                    lut_structure[25]  = 32'h0D14E3BC;
                    lut_structure[26]  = 32'h0CD9E83E;
                    lut_structure[27]  = 32'h0C9CE075;
                    lut_structure[28]  = 32'h0C5E353F;
                    lut_structure[29]  = 32'h0C1D7DBF;
                    lut_structure[30]  = 32'h0BDB22D0;
                    lut_structure[31]  = 32'h0B9652BD;
                    lut_structure[32]  = 32'h0B504816;
                    lut_structure[33]  = 32'h0B083126;
                    lut_structure[34]  = 32'h0ABEDFA4;
                    lut_structure[35]  = 32'h0A7381D7;
                    lut_structure[36]  = 32'h0A26809D;
                    lut_structure[37]  = 32'h09D7DBF4;
                    lut_structure[38]  = 32'h0987FCB9;
                    lut_structure[39]  = 32'h09367A0F;
                    lut_structure[40]  = 32'h08E3BCD3;
                    lut_structure[41]  = 32'h088F5C28;
                    lut_structure[42]  = 32'h0839C0EB;
                    lut_structure[43]  = 32'h07E2EB1C;
                    lut_structure[44]  = 32'h078ADAB9;
                    lut_structure[45]  = 32'h07318FC5;
                    lut_structure[46]  = 32'h06D77318;
                    lut_structure[47]  = 32'h067BB2FE;
                    lut_structure[48]  = 32'h061F8A09;
                    lut_structure[49]  = 32'h05C22680;
                    lut_structure[50]  = 32'h0563F141;
                    lut_structure[51]  = 32'h0504EA4A;
                    lut_structure[52]  = 32'h04A5119C;
                    lut_structure[53]  = 32'h04446738;
                    lut_structure[54]  = 32'h03E353F7;
                    lut_structure[55]  = 32'h03816F00;
                    lut_structure[56]  = 32'h031F212D;
                    lut_structure[57]  = 32'h02BC6A7E;
                    lut_structure[58]  = 32'h0258E219;
                    lut_structure[59]  = 32'h01F559B3;
                    lut_structure[60]  = 32'h01916872;
                    lut_structure[61]  = 32'h012D7731;
                    lut_structure[62]  = 32'h00C91D14;
                    lut_structure[63]  = 32'h00645A1C;
                    lut_structure[64]  = 32'h00000000;
                    lut_structure[65]  = 32'hFF9BA5E4;
                    lut_structure[66]  = 32'hFF36E2EC;
                    lut_structure[67]  = 32'hFED288CF;
                    lut_structure[68]  = 32'hFE6E978E;
                    lut_structure[69]  = 32'hFE0AA64D;
                    lut_structure[70]  = 32'hFDA71DE7;
                    lut_structure[71]  = 32'hFD439582;
                    lut_structure[72]  = 32'hFCE0DED3;
                    lut_structure[73]  = 32'hFC7E91FF;
                    lut_structure[74]  = 32'hFC1CAC09;
                    lut_structure[75]  = 32'hFBBB98C8;
                    lut_structure[76]  = 32'hFB5AEE64;
                    lut_structure[77]  = 32'hFAFB15B6;
                    lut_structure[78]  = 32'hFA9C0EBF;
                    lut_structure[79]  = 32'hFA3DD980;
                    lut_structure[80]  = 32'hF9E075F7;
                    lut_structure[81]  = 32'hF9844D02;
                    lut_structure[82]  = 32'hF9288CE8;
                    lut_structure[83]  = 32'hF8CE703B;
                    lut_structure[84]  = 32'hF8752547;
                    lut_structure[85]  = 32'hF81D14E4;
                    lut_structure[86]  = 32'hF7C63F15;
                    lut_structure[87]  = 32'hF770A3D8;
                    lut_structure[88]  = 32'hF71C432D;
                    lut_structure[89]  = 32'hF6C985F1;
                    lut_structure[90]  = 32'hF6780347;
                    lut_structure[91]  = 32'hF628240C;
                    lut_structure[92]  = 32'hF5D97F63;
                    lut_structure[93]  = 32'hF58C7E29;
                    lut_structure[94]  = 32'hF541205C;
                    lut_structure[95]  = 32'hF4F7CEDA;
                    lut_structure[96]  = 32'hF4AFB7EA;
                    lut_structure[97]  = 32'hF469AD43;
                    lut_structure[98]  = 32'hF424DD30;
                    lut_structure[99]  = 32'hF3E28241;
                    lut_structure[100] = 32'hF3A1CAC1;
                    lut_structure[101] = 32'hF3631F8B;
                    lut_structure[102] = 32'hF32617C2;
                    lut_structure[103] = 32'hF2EB1C44;
                    lut_structure[104] = 32'hF2B22D0F;
                    lut_structure[105] = 32'hF27B4A24;
                    lut_structure[106] = 32'hF246DC5E;
                    lut_structure[107] = 32'hF2141206;
                    lut_structure[108] = 32'hF1E3BCD4;
                    lut_structure[109] = 32'hF1B573EB;
                    lut_structure[110] = 32'hF189374C;
                    lut_structure[111] = 32'hF15F6FD3;
                    lut_structure[112] = 32'hF137B4A3;
                    lut_structure[113] = 32'hF1126E98;
                    lut_structure[114] = 32'hF0EF9DB3;
                    lut_structure[115] = 32'hF0CED917;
                    lut_structure[116] = 32'hF0B089A1;
                    lut_structure[117] = 32'hF0944674;
                    lut_structure[118] = 32'hF07AE148;
                    lut_structure[119] = 32'hF0638866;
                    lut_structure[120] = 32'hF04EA4A9;
                    lut_structure[121] = 32'hF03C3612;
                    lut_structure[122] = 32'hF02C3C9F;
                    lut_structure[123] = 32'hF01EB852;
                    lut_structure[124] = 32'hF013A92B;
                    lut_structure[125] = 32'hF00B0F28;
                    lut_structure[126] = 32'hF004EA4B;
                    lut_structure[127] = 32'hF0013A93;
                    lut_structure[128] = 32'hF0000000;
                    lut_structure[129] = 32'hF0013A93;
                    lut_structure[130] = 32'hF004EA4B;
                    lut_structure[131] = 32'hF00B0F28;
                    lut_structure[132] = 32'hF013A92B;
                    lut_structure[133] = 32'hF01EB852;
                    lut_structure[134] = 32'hF02C3C9F;
                    lut_structure[135] = 32'hF03C3612;
                    lut_structure[136] = 32'hF04EA4A9;
                    lut_structure[137] = 32'hF0638866;
                    lut_structure[138] = 32'hF07AE148;
                    lut_structure[139] = 32'hF0944674;
                    lut_structure[140] = 32'hF0B089A1;
                    lut_structure[141] = 32'hF0CED917;
                    lut_structure[142] = 32'hF0EF9DB3;
                    lut_structure[143] = 32'hF1126E98;
                    lut_structure[144] = 32'hF137B4A3;
                    lut_structure[145] = 32'hF15F6FD3;
                    lut_structure[146] = 32'hF189374C;
                    lut_structure[147] = 32'hF1B573EB;
                    lut_structure[148] = 32'hF1E3BCD4;
                    lut_structure[149] = 32'hF2141206;
                    lut_structure[150] = 32'hF246DC5E;
                    lut_structure[151] = 32'hF27B4A24;
                    lut_structure[152] = 32'hF2B22D0F;
                    lut_structure[153] = 32'hF2EB1C44;
                    lut_structure[154] = 32'hF32617C2;
                    lut_structure[155] = 32'hF3631F8B;
                    lut_structure[156] = 32'hF3A1CAC1;
                    lut_structure[157] = 32'hF3E28241;
                    lut_structure[158] = 32'hF424DD30;
                    lut_structure[159] = 32'hF469AD43;
                    lut_structure[160] = 32'hF4AFB7EA;
                    lut_structure[161] = 32'hF4F7CEDA;
                    lut_structure[162] = 32'hF541205C;
                    lut_structure[163] = 32'hF58C7E29;
                    lut_structure[164] = 32'hF5D97F63;
                    lut_structure[165] = 32'hF628240C;
                    lut_structure[166] = 32'hF6780347;
                    lut_structure[167] = 32'hF6C985F1;
                    lut_structure[168] = 32'hF71C432D;
                    lut_structure[169] = 32'hF770A3D8;
                    lut_structure[170] = 32'hF7C63F15;
                    lut_structure[171] = 32'hF81D14E4;
                    lut_structure[172] = 32'hF8752547;
                    lut_structure[173] = 32'hF8CE703B;
                    lut_structure[174] = 32'hF9288CE8;
                    lut_structure[175] = 32'hF9844D02;
                    lut_structure[176] = 32'hF9E075F7;
                    lut_structure[177] = 32'hFA3DD980;
                    lut_structure[178] = 32'hFA9C0EBF;
                    lut_structure[179] = 32'hFAFB15B6;
                    lut_structure[180] = 32'hFB5AEE64;
                    lut_structure[181] = 32'hFBBB98C8;
                    lut_structure[182] = 32'hFC1CAC09;
                    lut_structure[183] = 32'hFC7E91FF;
                    lut_structure[184] = 32'hFCE0DED3;
                    lut_structure[185] = 32'hFD439582;
                    lut_structure[186] = 32'hFDA71DE7;
                    lut_structure[187] = 32'hFE0AA64D;
                    lut_structure[188] = 32'hFE6E978E;
                    lut_structure[189] = 32'hFED288CF;
                    lut_structure[190] = 32'hFF36E2EC;
                    lut_structure[191] = 32'hFF9BA5E4;
                    lut_structure[192] = 32'h00000000;
                    lut_structure[193] = 32'h00645A1C;
                    lut_structure[194] = 32'h00C91D14;
                    lut_structure[195] = 32'h012D7731;
                    lut_structure[196] = 32'h01916872;
                    lut_structure[197] = 32'h01F559B3;
                    lut_structure[198] = 32'h0258E219;
                    lut_structure[199] = 32'h02BC6A7E;
                    lut_structure[200] = 32'h031F212D;
                    lut_structure[201] = 32'h03816F00;
                    lut_structure[202] = 32'h03E353F7;
                    lut_structure[203] = 32'h04446738;
                    lut_structure[204] = 32'h04A5119C;
                    lut_structure[205] = 32'h0504EA4A;
                    lut_structure[206] = 32'h0563F141;
                    lut_structure[207] = 32'h05C22680;
                    lut_structure[208] = 32'h061F8A09;
                    lut_structure[209] = 32'h067BB2FE;
                    lut_structure[210] = 32'h06D77318;
                    lut_structure[211] = 32'h07318FC5;
                    lut_structure[212] = 32'h078ADAB9;
                    lut_structure[213] = 32'h07E2EB1C;
                    lut_structure[214] = 32'h0839C0EB;
                    lut_structure[215] = 32'h088F5C28;
                    lut_structure[216] = 32'h08E3BCD3;
                    lut_structure[217] = 32'h09367A0F;
                    lut_structure[218] = 32'h0987FCB9;
                    lut_structure[219] = 32'h09D7DBF4;
                    lut_structure[220] = 32'h0A26809D;
                    lut_structure[221] = 32'h0A7381D7;
                    lut_structure[222] = 32'h0ABEDFA4;
                    lut_structure[223] = 32'h0B083126;
                    lut_structure[224] = 32'h0B504816;
                    lut_structure[225] = 32'h0B9652BD;
                    lut_structure[226] = 32'h0BDB22D0;
                    lut_structure[227] = 32'h0C1D7DBF;
                    lut_structure[228] = 32'h0C5E353F;
                    lut_structure[229] = 32'h0C9CE075;
                    lut_structure[230] = 32'h0CD9E83E;
                    lut_structure[231] = 32'h0D14E3BC;
                    lut_structure[232] = 32'h0D4DD2F1;
                    lut_structure[233] = 32'h0D84B5DC;
                    lut_structure[234] = 32'h0DB923A2;
                    lut_structure[235] = 32'h0DEBEDFA;
                    lut_structure[236] = 32'h0E1C432C;
                    lut_structure[237] = 32'h0E4A8C15;
                    lut_structure[238] = 32'h0E76C8B4;
                    lut_structure[239] = 32'h0EA0902D;
                    lut_structure[240] = 32'h0EC84B5D;
                    lut_structure[241] = 32'h0EED9168;
                    lut_structure[242] = 32'h0F10624D;
                    lut_structure[243] = 32'h0F3126E9;
                    lut_structure[244] = 32'h0F4F765F;
                    lut_structure[245] = 32'h0F6BB98C;
                    lut_structure[246] = 32'h0F851EB8;
                    lut_structure[247] = 32'h0F9C779A;
                    lut_structure[248] = 32'h0FB15B57;
                    lut_structure[249] = 32'h0FC3C9EE;
                    lut_structure[250] = 32'h0FD3C361;
                    lut_structure[251] = 32'h0FE147AE;
                    lut_structure[252] = 32'h0FEC56D5;
                    lut_structure[253] = 32'h0FF4F0D8;
                    lut_structure[254] = 32'h0FFB15B5;
                    lut_structure[255] = 32'h0FFEC56D;


                end
                //trian
                else if(TXT_FILE == 3) begin 
                    lut_structure[0]   = 32'h00000000;
                    lut_structure[1]   = 32'h003FE5C9;
                    lut_structure[2]   = 32'h007FCB92;
                    lut_structure[3]   = 32'h00C01A36;
                    lut_structure[4]   = 32'h01000000;
                    lut_structure[5]   = 32'h013FE5C9;
                    lut_structure[6]   = 32'h0180346D;
                    lut_structure[7]   = 32'h01C01A36;
                    lut_structure[8]   = 32'h02000000;
                    lut_structure[9]   = 32'h023FE5C9;
                    lut_structure[10]  = 32'h027FCB92;
                    lut_structure[11]  = 32'h02C01A36;
                    lut_structure[12]  = 32'h03000000;
                    lut_structure[13]  = 32'h033FE5C9;
                    lut_structure[14]  = 32'h0380346D;
                    lut_structure[15]  = 32'h03C01A36;
                    lut_structure[16]  = 32'h04000000;
                    lut_structure[17]  = 32'h043FE5C9;
                    lut_structure[18]  = 32'h047FCB92;
                    lut_structure[19]  = 32'h04C01A36;
                    lut_structure[20]  = 32'h05000000;
                    lut_structure[21]  = 32'h053FE5C9;
                    lut_structure[22]  = 32'h0580346D;
                    lut_structure[23]  = 32'h05C01A36;
                    lut_structure[24]  = 32'h06000000;
                    lut_structure[25]  = 32'h063FE5C9;
                    lut_structure[26]  = 32'h067FCB92;
                    lut_structure[27]  = 32'h06C01A36;
                    lut_structure[28]  = 32'h07000000;
                    lut_structure[29]  = 32'h073FE5C9;
                    lut_structure[30]  = 32'h0780346D;
                    lut_structure[31]  = 32'h07C01A36;
                    lut_structure[32]  = 32'h08000000;
                    lut_structure[33]  = 32'h083FE5C9;
                    lut_structure[34]  = 32'h087FCB92;
                    lut_structure[35]  = 32'h08C01A36;
                    lut_structure[36]  = 32'h09000000;
                    lut_structure[37]  = 32'h093FE5C9;
                    lut_structure[38]  = 32'h0980346D;
                    lut_structure[39]  = 32'h09C01A36;
                    lut_structure[40]  = 32'h0A000000;
                    lut_structure[41]  = 32'h0A3FE5C9;
                    lut_structure[42]  = 32'h0A7FCB92;
                    lut_structure[43]  = 32'h0AC01A36;
                    lut_structure[44]  = 32'h0B000000;
                    lut_structure[45]  = 32'h0B3FE5C9;
                    lut_structure[46]  = 32'h0B80346D;
                    lut_structure[47]  = 32'h0BC01A36;
                    lut_structure[48]  = 32'h0C000000;
                    lut_structure[49]  = 32'h0C3FE5C9;
                    lut_structure[50]  = 32'h0C7FCB92;
                    lut_structure[51]  = 32'h0CC01A36;
                    lut_structure[52]  = 32'h0D000000;
                    lut_structure[53]  = 32'h0D3FE5C9;
                    lut_structure[54]  = 32'h0D80346D;
                    lut_structure[55]  = 32'h0DC01A36;
                    lut_structure[56]  = 32'h0E000000;
                    lut_structure[57]  = 32'h0E3FE5C9;
                    lut_structure[58]  = 32'h0E3FE5C9;
                    lut_structure[59]  = 32'h0EC01A36;
                    lut_structure[60]  = 32'h0F000000;
                    lut_structure[61]  = 32'h0F3FE5C9;
                    lut_structure[62]  = 32'h0F80346D;
                    lut_structure[63]  = 32'h0FC01A36;
                    lut_structure[64]  = 32'h10000000;
                    lut_structure[65]  = 32'h0FC01A36;
                    lut_structure[66]  = 32'h0F80346D;
                    lut_structure[67]  = 32'h0F3FE5C9;
                    lut_structure[68]  = 32'h0F000000;
                    lut_structure[69]  = 32'h0EC01A36;
                    lut_structure[70]  = 32'h0E7FCB92;
                    lut_structure[71]  = 32'h0E3FE5C9;
                    lut_structure[72]  = 32'h0E000000;
                    lut_structure[73]  = 32'h0DC01A36;
                    lut_structure[74]  = 32'h0D80346D;
                    lut_structure[75]  = 32'h0D3FE5C9;
                    lut_structure[76]  = 32'h0D000000;
                    lut_structure[77]  = 32'h0CC01A36;
                    lut_structure[78]  = 32'h0C7FCB92;
                    lut_structure[79]  = 32'h0C3FE5C9;
                    lut_structure[80]  = 32'h0C000000;
                    lut_structure[81]  = 32'h0BC01A36;
                    lut_structure[82]  = 32'h0B80346D;
                    lut_structure[83]  = 32'h0B3FE5C9;
                    lut_structure[84]  = 32'h0B000000;
                    lut_structure[85]  = 32'h0AC01A36;
                    lut_structure[86]  = 32'h0A7BCB92;
                    lut_structure[87]  = 32'h0A3FE5C9;
                    lut_structure[88]  = 32'h0A000000;
                    lut_structure[89]  = 32'h09C01A36;
                    lut_structure[90]  = 32'h0980346D;
                    lut_structure[91]  = 32'h093FE5C9;
                    lut_structure[92]  = 32'h09000000;
                    lut_structure[93]  = 32'h08C01A36;
                    lut_structure[94]  = 32'h087FCB92;
                    lut_structure[95]  = 32'h083FE5C9;
                    lut_structure[96]  = 32'h08000000;
                    lut_structure[97]  = 32'h07C01A36;
                    lut_structure[98]  = 32'h0780346D;
                    lut_structure[99]  = 32'h073FE5C9;
                    lut_structure[100] = 32'h07000000;
                    lut_structure[101] = 32'h06C01A36;
                    lut_structure[102] = 32'h067FCB92;
                    lut_structure[103] = 32'h063FE5C9;
                    lut_structure[104] = 32'h06000000;
                    lut_structure[105] = 32'h05C01A36;
                    lut_structure[106] = 32'h0580346D;
                    lut_structure[107] = 32'h053FE5C9;
                    lut_structure[108] = 32'h05000000;
                    lut_structure[109] = 32'h04C01A36;
                    lut_structure[110] = 32'h047FCB92;
                    lut_structure[111] = 32'h043FE5C9;
                    lut_structure[112] = 32'h04000000;
                    lut_structure[113] = 32'h03C01A36;
                    lut_structure[114] = 32'h0380346D;
                    lut_structure[115] = 32'h033FE5C9;
                    lut_structure[116] = 32'h03000000;
                    lut_structure[117] = 32'h02C01A36;
                    lut_structure[118] = 32'h027FCB92;
                    lut_structure[119] = 32'h023FE5C9;
                    lut_structure[120] = 32'h02000000;
                    lut_structure[121] = 32'h01C01A36;
                    lut_structure[122] = 32'h0180346D;
                    lut_structure[123] = 32'h013FE5C9;
                    lut_structure[124] = 32'h01000000;
                    lut_structure[125] = 32'h00C01A36;
                    lut_structure[126] = 32'h007FCB92;
                    lut_structure[127] = 32'h003FE5C9;
                    lut_structure[128] = 32'h00000000;
                    lut_structure[129] = 32'hFFC01A37;
                    lut_structure[130] = 32'hFF80346E;
                    lut_structure[131] = 32'hFF3FE5CA;
                    lut_structure[132] = 32'hFF000000;
                    lut_structure[133] = 32'hFEC01A37;
                    lut_structure[134] = 32'hFE7FCB93;
                    lut_structure[135] = 32'hFE3FE5CA;
                    lut_structure[136] = 32'hFE000000;
                    lut_structure[137] = 32'hFDC01A37;
                    lut_structure[138] = 32'hFD80346E;
                    lut_structure[139] = 32'hFD3FE5CA;
                    lut_structure[140] = 32'hFD000000;
                    lut_structure[141] = 32'hFCC01A37;
                    lut_structure[142] = 32'hFC7FCB93;
                    lut_structure[143] = 32'hFC3FE5CA;
                    lut_structure[144] = 32'hFC000000;
                    lut_structure[145] = 32'hFBC01A37;
                    lut_structure[146] = 32'hFB80346E;
                    lut_structure[147] = 32'hFB3FE5CA;
                    lut_structure[148] = 32'hFB000000;
                    lut_structure[149] = 32'hFAC01A37;
                    lut_structure[150] = 32'hFA7BCB93;
                    lut_structure[151] = 32'hFA3FE5CA;
                    lut_structure[152] = 32'hFA000000;
                    lut_structure[153] = 32'hF9C01A37;
                    lut_structure[154] = 32'hF980346E;
                    lut_structure[155] = 32'hF93FE5CA;
                    lut_structure[156] = 32'hF9000000;
                    lut_structure[157] = 32'hF8C01A37;
                    lut_structure[158] = 32'hF87FCB93;
                    lut_structure[159] = 32'hF83FE5CA;
                    lut_structure[160] = 32'hF8000000;
                    lut_structure[161] = 32'hF7C01A37;
                    lut_structure[162] = 32'hF780346E;
                    lut_structure[163] = 32'hF73FE5CA;
                    lut_structure[164] = 32'hF7000000;
                    lut_structure[165] = 32'hF6C01A37;
                    lut_structure[166] = 32'hF67FCB93;
                    lut_structure[167] = 32'hF63FE5CA;
                    lut_structure[168] = 32'hF6000000;
                    lut_structure[169] = 32'hF5C01A37;
                    lut_structure[170] = 32'hF580346E;
                    lut_structure[171] = 32'hF53FE5CA;
                    lut_structure[172] = 32'hF5000000;
                    lut_structure[173] = 32'hF4C01A37;
                    lut_structure[174] = 32'hF47FCB93;
                    lut_structure[175] = 32'hF43FE5CA;
                    lut_structure[176] = 32'hF4000000;
                    lut_structure[177] = 32'hF3C01A37;
                    lut_structure[178] = 32'hF380346E;
                    lut_structure[179] = 32'hF33FE5CA;
                    lut_structure[180] = 32'hF3000000;
                    lut_structure[181] = 32'hF2C01A37;
                    lut_structure[182] = 32'hF27FCB93;
                    lut_structure[183] = 32'hF23FE5CA;
                    lut_structure[184] = 32'hF2000000;
                    lut_structure[185] = 32'hF1C01A37;
                    lut_structure[186] = 32'hF180346E;
                    lut_structure[187] = 32'hF13FE5CA;
                    lut_structure[188] = 32'hF1000000;
                    lut_structure[189] = 32'hF0C01A37;
                    lut_structure[190] = 32'hF07FCB93;
                    lut_structure[191] = 32'hF03FE5CA;
                    lut_structure[192] = 32'hF0000000;
                    lut_structure[193] = 32'hF03FE5CA;
                    lut_structure[194] = 32'hF07FCB93;
                    lut_structure[195] = 32'hF0C01A37;
                    lut_structure[196] = 32'hF1000000;
                    lut_structure[197] = 32'hF13FE5CA;
                    lut_structure[198] = 32'hF180346E;
                    lut_structure[199] = 32'hF1C01A37;
                    lut_structure[200] = 32'hF2000000;
                    lut_structure[201] = 32'hF23FE5CA;
                    lut_structure[202] = 32'hF27FCB93;
                    lut_structure[203] = 32'hF2C01A37;
                    lut_structure[204] = 32'hF3000000;
                    lut_structure[205] = 32'hF33FE5CA;
                    lut_structure[206] = 32'hF380346E;
                    lut_structure[207] = 32'hF3C01A37;
                    lut_structure[208] = 32'hF4000000;
                    lut_structure[209] = 32'hF43FE5CA;
                    lut_structure[210] = 32'hF47FCB93;
                    lut_structure[211] = 32'hF4C01A37;
                    lut_structure[212] = 32'hF5000000;
                    lut_structure[213] = 32'hF53FE5CA;
                    lut_structure[214] = 32'hF580346E;
                    lut_structure[215] = 32'hF5C01A37;
                    lut_structure[216] = 32'hF6000000;
                    lut_structure[217] = 32'hF63FE5CA;
                    lut_structure[218] = 32'hF67FCB93;
                    lut_structure[219] = 32'hF6C01A37;
                    lut_structure[220] = 32'hF7000000;
                    lut_structure[221] = 32'hF73FE5CA;
                    lut_structure[222] = 32'hF780346E;
                    lut_structure[223] = 32'hF7C01A37;
                    lut_structure[224] = 32'hF8000000;
                    lut_structure[225] = 32'hF83FE5CA;
                    lut_structure[226] = 32'hF87FCB93;
                    lut_structure[227] = 32'hF8C01A37;
                    lut_structure[228] = 32'hF9000000;
                    lut_structure[229] = 32'hF93FE5CA;
                    lut_structure[230] = 32'hF980346E;
                    lut_structure[231] = 32'hF9C01A37;
                    lut_structure[232] = 32'hFA000000;
                    lut_structure[233] = 32'hFA3FE5CA;
                    lut_structure[234] = 32'hFA7FCB93;
                    lut_structure[235] = 32'hFAC01A37;
                    lut_structure[236] = 32'hFB000000;
                    lut_structure[237] = 32'hFB3FE5CA;
                    lut_structure[238] = 32'hFB80346E;
                    lut_structure[239] = 32'hFBC01A37;
                    lut_structure[240] = 32'hFC000000;
                    lut_structure[241] = 32'hFC3FE5CA;
                    lut_structure[242] = 32'hFC7FCB93;
                    lut_structure[243] = 32'hFCC01A37;
                    lut_structure[244] = 32'hFD000000;
                    lut_structure[245] = 32'hFD3FE5CA;
                    lut_structure[246] = 32'hFD80346E;
                    lut_structure[247] = 32'hFDC01A37;
                    lut_structure[248] = 32'hFE000000;
                    lut_structure[249] = 32'hFE3FE5CA;
                    lut_structure[250] = 32'hFE7FCB93;
                    lut_structure[251] = 32'hFEC01A37;
                    lut_structure[252] = 32'hFF000000;
                    lut_structure[253] = 32'hFF3FE5CA;
                    lut_structure[254] = 32'hFF80346E;
                    lut_structure[255] = 32'hFFC01A37;
                end                          
                //squa
                else if(TXT_FILE == 4) begin 
                    lut_structure[0]   = 32'h10000000;
                    lut_structure[1]   = 32'h10000000;
                    lut_structure[2]   = 32'h10000000;
                    lut_structure[3]   = 32'h10000000;
                    lut_structure[4]   = 32'h10000000;
                    lut_structure[5]   = 32'h10000000;
                    lut_structure[6]   = 32'h10000000;
                    lut_structure[7]   = 32'h10000000;
                    lut_structure[8]   = 32'h10000000;
                    lut_structure[9]   = 32'h10000000;
                    lut_structure[10]  = 32'h10000000;
                    lut_structure[11]  = 32'h10000000;
                    lut_structure[12]  = 32'h10000000;
                    lut_structure[13]  = 32'h10000000;
                    lut_structure[14]  = 32'h10000000;
                    lut_structure[15]  = 32'h10000000;
                    lut_structure[16]  = 32'h10000000;
                    lut_structure[17]  = 32'h10000000;
                    lut_structure[18]  = 32'h10000000;
                    lut_structure[19]  = 32'h10000000;
                    lut_structure[20]  = 32'h10000000;
                    lut_structure[21]  = 32'h10000000;
                    lut_structure[22]  = 32'h10000000;
                    lut_structure[23]  = 32'h10000000;
                    lut_structure[24]  = 32'h10000000;
                    lut_structure[25]  = 32'h10000000;
                    lut_structure[26]  = 32'h10000000;
                    lut_structure[27]  = 32'h10000000;
                    lut_structure[28]  = 32'h10000000;
                    lut_structure[29]  = 32'h10000000;
                    lut_structure[30]  = 32'h10000000;
                    lut_structure[31]  = 32'h10000000;
                    lut_structure[32]  = 32'h10000000;
                    lut_structure[33]  = 32'h10000000;
                    lut_structure[34]  = 32'h10000000;
                    lut_structure[35]  = 32'h10000000;
                    lut_structure[36]  = 32'h10000000;
                    lut_structure[37]  = 32'h10000000;
                    lut_structure[38]  = 32'h10000000;
                    lut_structure[39]  = 32'h10000000;
                    lut_structure[40]  = 32'h10000000;
                    lut_structure[41]  = 32'h10000000;
                    lut_structure[42]  = 32'h10000000;
                    lut_structure[43]  = 32'h10000000;
                    lut_structure[44]  = 32'h10000000;
                    lut_structure[45]  = 32'h10000000;
                    lut_structure[46]  = 32'h10000000;
                    lut_structure[47]  = 32'h10000000;
                    lut_structure[48]  = 32'h10000000;
                    lut_structure[49]  = 32'h10000000;
                    lut_structure[50]  = 32'h10000000;
                    lut_structure[51]  = 32'h10000000;
                    lut_structure[52]  = 32'h10000000;
                    lut_structure[53]  = 32'h10000000;
                    lut_structure[54]  = 32'h10000000;
                    lut_structure[55]  = 32'h10000000;
                    lut_structure[56]  = 32'h10000000;
                    lut_structure[57]  = 32'h10000000;
                    lut_structure[58]  = 32'h10000000;
                    lut_structure[59]  = 32'h10000000;
                    lut_structure[60]  = 32'h10000000;
                    lut_structure[61]  = 32'h10000000;
                    lut_structure[62]  = 32'h10000000;
                    lut_structure[63]  = 32'h10000000;
                    lut_structure[64]  = 32'h10000000;
                    lut_structure[65]  = 32'h10000000;
                    lut_structure[66]  = 32'h10000000;
                    lut_structure[67]  = 32'h10000000;
                    lut_structure[68]  = 32'h10000000;
                    lut_structure[69]  = 32'h10000000;
                    lut_structure[70]  = 32'h10000000;
                    lut_structure[71]  = 32'h10000000;
                    lut_structure[72]  = 32'h10000000;
                    lut_structure[73]  = 32'h10000000;
                    lut_structure[74]  = 32'h10000000;
                    lut_structure[75]  = 32'h10000000;
                    lut_structure[76]  = 32'h10000000;
                    lut_structure[77]  = 32'h10000000;
                    lut_structure[78]  = 32'h10000000;
                    lut_structure[79]  = 32'h10000000;
                    lut_structure[80]  = 32'h10000000;
                    lut_structure[81]  = 32'h10000000;
                    lut_structure[82]  = 32'h10000000;
                    lut_structure[83]  = 32'h10000000;
                    lut_structure[84]  = 32'h10000000;
                    lut_structure[85]  = 32'h10000000;
                    lut_structure[86]  = 32'h10000000;
                    lut_structure[87]  = 32'h10000000;
                    lut_structure[88]  = 32'h10000000;
                    lut_structure[89]  = 32'h10000000;
                    lut_structure[90]  = 32'h10000000;
                    lut_structure[91]  = 32'h10000000;
                    lut_structure[92]  = 32'h10000000;
                    lut_structure[93]  = 32'h10000000;
                    lut_structure[94]  = 32'h10000000;
                    lut_structure[95]  = 32'h10000000;
                    lut_structure[96]  = 32'h10000000;
                    lut_structure[97]  = 32'h10000000;
                    lut_structure[98]  = 32'h10000000;
                    lut_structure[99]  = 32'h10000000;
                    lut_structure[100] = 32'h10000000;
                    lut_structure[101] = 32'h10000000;
                    lut_structure[102] = 32'h10000000;
                    lut_structure[103] = 32'h10000000;
                    lut_structure[104] = 32'h10000000;
                    lut_structure[105] = 32'h10000000;
                    lut_structure[106] = 32'h10000000;
                    lut_structure[107] = 32'h10000000;
                    lut_structure[108] = 32'h10000000;
                    lut_structure[109] = 32'h10000000;
                    lut_structure[110] = 32'h10000000;
                    lut_structure[111] = 32'h10000000;
                    lut_structure[112] = 32'h10000000;
                    lut_structure[113] = 32'h10000000;
                    lut_structure[114] = 32'h10000000;
                    lut_structure[115] = 32'h10000000;
                    lut_structure[116] = 32'h10000000;
                    lut_structure[117] = 32'h10000000;
                    lut_structure[118] = 32'h10000000;
                    lut_structure[119] = 32'h10000000;
                    lut_structure[120] = 32'h10000000;
                    lut_structure[121] = 32'h10000000;
                    lut_structure[122] = 32'h10000000;
                    lut_structure[123] = 32'h10000000;
                    lut_structure[124] = 32'h10000000;
                    lut_structure[125] = 32'h10000000;
                    lut_structure[126] = 32'h10000000;
                    lut_structure[127] = 32'h10000000;
                    lut_structure[128] = 32'hF0000000;
                    lut_structure[129] = 32'hF0000000;
                    lut_structure[130] = 32'hF0000000;
                    lut_structure[131] = 32'hF0000000;
                    lut_structure[132] = 32'hF0000000;
                    lut_structure[133] = 32'hF0000000;
                    lut_structure[134] = 32'hF0000000;
                    lut_structure[135] = 32'hF0000000;
                    lut_structure[136] = 32'hF0000000;
                    lut_structure[137] = 32'hF0000000;
                    lut_structure[138] = 32'hF0000000;
                    lut_structure[139] = 32'hF0000000;
                    lut_structure[140] = 32'hF0000000;
                    lut_structure[141] = 32'hF0000000;
                    lut_structure[142] = 32'hF0000000;
                    lut_structure[143] = 32'hF0000000;
                    lut_structure[144] = 32'hF0000000;
                    lut_structure[145] = 32'hF0000000;
                    lut_structure[146] = 32'hF0000000;
                    lut_structure[147] = 32'hF0000000;
                    lut_structure[148] = 32'hF0000000;
                    lut_structure[149] = 32'hF0000000;
                    lut_structure[150] = 32'hF0000000;
                    lut_structure[151] = 32'hF0000000;
                    lut_structure[152] = 32'hF0000000;
                    lut_structure[153] = 32'hF0000000;
                    lut_structure[154] = 32'hF0000000;
                    lut_structure[155] = 32'hF0000000;
                    lut_structure[156] = 32'hF0000000;
                    lut_structure[157] = 32'hF0000000;
                    lut_structure[158] = 32'hF0000000;
                    lut_structure[159] = 32'hF0000000;
                    lut_structure[160] = 32'hF0000000;
                    lut_structure[161] = 32'hF0000000;
                    lut_structure[162] = 32'hF0000000;
                    lut_structure[163] = 32'hF0000000;
                    lut_structure[164] = 32'hF0000000;
                    lut_structure[165] = 32'hF0000000;
                    lut_structure[166] = 32'hF0000000;
                    lut_structure[167] = 32'hF0000000;
                    lut_structure[168] = 32'hF0000000;
                    lut_structure[169] = 32'hF0000000;
                    lut_structure[170] = 32'hF0000000;
                    lut_structure[171] = 32'hF0000000;
                    lut_structure[172] = 32'hF0000000;
                    lut_structure[173] = 32'hF0000000;
                    lut_structure[174] = 32'hF0000000;
                    lut_structure[175] = 32'hF0000000;
                    lut_structure[176] = 32'hF0000000;
                    lut_structure[177] = 32'hF0000000;
                    lut_structure[178] = 32'hF0000000;
                    lut_structure[179] = 32'hF0000000;
                    lut_structure[180] = 32'hF0000000;
                    lut_structure[181] = 32'hF0000000;
                    lut_structure[182] = 32'hF0000000;
                    lut_structure[183] = 32'hF0000000;
                    lut_structure[184] = 32'hF0000000;
                    lut_structure[185] = 32'hF0000000;
                    lut_structure[186] = 32'hF0000000;
                    lut_structure[187] = 32'hF0000000;
                    lut_structure[188] = 32'hF0000000;
                    lut_structure[189] = 32'hF0000000;
                    lut_structure[190] = 32'hF0000000;
                    lut_structure[191] = 32'hF0000000;
                    lut_structure[192] = 32'hF0000000;
                    lut_structure[193] = 32'hF0000000;
                    lut_structure[194] = 32'hF0000000;
                    lut_structure[195] = 32'hF0000000;
                    lut_structure[196] = 32'hF0000000;
                    lut_structure[197] = 32'hF0000000;
                    lut_structure[198] = 32'hF0000000;
                    lut_structure[199] = 32'hF0000000;
                    lut_structure[200] = 32'hF0000000;
                    lut_structure[201] = 32'hF0000000;
                    lut_structure[202] = 32'hF0000000;
                    lut_structure[203] = 32'hF0000000;
                    lut_structure[204] = 32'hF0000000;
                    lut_structure[205] = 32'hF0000000;
                    lut_structure[206] = 32'hF0000000;
                    lut_structure[207] = 32'hF0000000;
                    lut_structure[208] = 32'hF0000000;
                    lut_structure[209] = 32'hF0000000;
                    lut_structure[210] = 32'hF0000000;
                    lut_structure[211] = 32'hF0000000;
                    lut_structure[212] = 32'hF0000000;
                    lut_structure[213] = 32'hF0000000;
                    lut_structure[214] = 32'hF0000000;
                    lut_structure[215] = 32'hF0000000;
                    lut_structure[216] = 32'hF0000000;
                    lut_structure[217] = 32'hF0000000;
                    lut_structure[218] = 32'hF0000000;
                    lut_structure[219] = 32'hF0000000;
                    lut_structure[220] = 32'hF0000000;
                    lut_structure[221] = 32'hF0000000;
                    lut_structure[222] = 32'hF0000000;
                    lut_structure[223] = 32'hF0000000;
                    lut_structure[224] = 32'hF0000000;
                    lut_structure[225] = 32'hF0000000;
                    lut_structure[226] = 32'hF0000000;
                    lut_structure[227] = 32'hF0000000;
                    lut_structure[228] = 32'hF0000000;
                    lut_structure[229] = 32'hF0000000;
                    lut_structure[230] = 32'hF0000000;
                    lut_structure[231] = 32'hF0000000;
                    lut_structure[232] = 32'hF0000000;
                    lut_structure[233] = 32'hF0000000;
                    lut_structure[234] = 32'hF0000000;
                    lut_structure[235] = 32'hF0000000;
                    lut_structure[236] = 32'hF0000000;
                    lut_structure[237] = 32'hF0000000;
                    lut_structure[238] = 32'hF0000000;
                    lut_structure[239] = 32'hF0000000;
                    lut_structure[240] = 32'hF0000000;
                    lut_structure[241] = 32'hF0000000;
                    lut_structure[242] = 32'hF0000000;
                    lut_structure[243] = 32'hF0000000;
                    lut_structure[244] = 32'hF0000000;
                    lut_structure[245] = 32'hF0000000;
                    lut_structure[246] = 32'hF0000000;
                    lut_structure[247] = 32'hF0000000;
                    lut_structure[248] = 32'hF0000000;
                    lut_structure[249] = 32'hF0000000;
                    lut_structure[250] = 32'hF0000000;
                    lut_structure[251] = 32'hF0000000;
                    lut_structure[252] = 32'hF0000000;
                    lut_structure[253] = 32'hF0000000;
                    lut_structure[254] = 32'hF0000000;
                    lut_structure[255] = 32'hF0000000;
                end
end
*/
//read operation
always_ff @ (posedge clk) begin	
		read_data_o <= lut_structure[read_addr_i];		
end

endmodule

